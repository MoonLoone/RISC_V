package tb_constants;
localparam int MEMORY_SIZE = 32;
localparam time CLK_PERIOD = 10;
localparam logic[31:0] SIM_STOP_PC = 24;
localparam int MEM_CHECK_ADDR = 64;
localparam logic[31:0] EXPECTED_RESULT = 49;
endpackage
